module apb_decoder (



);



endmodule

/* APB Header file */
`define TOTAL_SLAVE 16

module top_apb (
input clk,
output pclk,
output pwdata
);

endmodule

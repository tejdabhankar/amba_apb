module apb_decoder (
	input clk,
	input f_empty,
	output rd_en,
	input fifo_data
	
);



endmodule
